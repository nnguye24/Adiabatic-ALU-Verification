`include "adder/custom_tranif.sv"
`include "adder/inv.sv"
`include "adder/inv_fo16.sv"
`include "adder/and2b.sv"
`include "adder/black_cell2b.sv"
`include "adder/black_cell_inv2b.sv"
`include "adder/gray_cell2b.sv"
`include "adder/gray_cell_inv2b.sv"
`include "adder/adder.sv"
`include "adder/bennettClock.sv"

module adder_b (
    input wire [15:0] a,      // 16-bit input
    input wire [15:0] b,      // 16-bit input
    input wire cin,
    input wire clk,      
    input wire reset,          
    output wire [15:0] out,   // Changed to wire
    output wire cout,
    output wire calculation_done,  // Signal for when result is valid
    output wire [7:0] clkp_out,    // Outputs for monitoring clock signals
    output wire [7:0] clkn_out,
    output wire [15:0] propagate,  // Expose propagate signals for verification
    output wire [15:0] generate_   // Expose generate signals for verification (note trailing underscore to avoid keyword)
);
    // Power supplies
    supply1 vdd;             
    supply0 vss;

    // Bennett clock signals
    wire instFlag;
    wire [7:0] clkneg;
    wire [7:0] clkpos;

    // Connect monitor outputs to internal clock signals
    assign clkp_out = clkpos;
    assign clkn_out = clkneg;

    // Bennett clock generator
    bennett_clock #(
        .WIDTH(8)  
    ) bennett_gen (
        .clk(clk),
        .reset(reset),
        .instFlag(instFlag),
        .clkn(clkneg),
        .clkp(clkpos)
    );

    wire [15:0] internal_p1;
    
    // Adder instance with individual port connections
    adder adder_inst ( 
        a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8],
        a[9], a[10], a[11], a[12], a[13], a[14], a[15], 
        b[0], b[1], b[2], b[3], b[4], b[5], b[6], b[7], b[8], 
        b[9], b[10], b[11], b[12], b[13], b[14], b[15], 
        cin, clkneg[0], clkneg[1], clkneg[2], clkneg[3], clkneg[4], 
        clkneg[5], clkneg[6], clkneg[7], clkpos[0], clkpos[1], 
        clkpos[2], clkpos[3], clkpos[4], clkpos[5], clkpos[6],
        clkpos[7], cout, out[0], out[1], out[2], out[3], out[4], 
        out[5], out[6], out[7], out[8], out[9], out[10], out[11], 
        out[12], out[13], out[14], out[15], vdd, vss
    );
    
    // Assign propagate and generate outputs
    // In this design, propagate signals are p = a XOR b
    // Generate signals are g = a AND b
    // We'll recreate them here since we can't directly access internal signals
    assign propagate = a ^ b;  // Propagate = a XOR b
    assign generate_ = a & b;  // Generate = a AND b
    
    // Signal to indicate when calculation is complete
    assign calculation_done = instFlag;
    
endmodule