package adder_pkg;
	import uvm_pkg::*;

	`include "adder_sequencer.sv"
	`include "adder_monitor.sv"
	`include "adder_driver.sv"
	`include "adder_agent.sv"
	`include "adder_scoreboard.sv"
	`include "adder_config.sv"
	`include "adder_env.sv"
	`include "adder_test.sv"
endpackage: adder_pkg